//
//File: json_object_test.svh
//Device: 
//Author: zhouchuanrui@foxmail.com
//Created:  2021/2/28 22:12:14
//Description: object test for json
//Revisions: 
//2021/2/28 22:12:24: created
//

