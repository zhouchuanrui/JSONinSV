//
//File: json_macros.svh
//Device: 
//Author: zhouchuanrui@foxmail.com
//Created:  2021/1/26 7:30:57
//Description: Macros for JSON lib
//Revisions: 
//2021/1/26 7:31:43: created
//

`define JSON_LOG()
`define JSON_WARN()
`define JSON_ERROR()
`define JSON_FATAL()

