//
//File: json_literal_test.svh
//Device: 
//Author: zhouchuanrui@foxmail.com
//Created:  2021/2/20 20:54:27
//Description: literal test for json
//Revisions: 
//2021/2/20 20:54:44: created
//

class json_literal_test extends TestPrototype;
    `__register(json_literal_test)

    task test();
        $display("Start JSON literal test..");
    endtask

endclass: json_literal_test

