//
//File: test_pkg.sv
//Device: 
//Created:  2017-4-18 22:55:14
//Description: test package
//Revisions: 
//2017-4-18 22:55:25: created
//

package test_pkg;
    `include "json_macros.svh"
    import json_pkg::JSONValue;

    `include "TestFactory.svh"
    `include "TestUtils.svh"
    `include "json_literal_test.svh"
    `include "json_string_test.svh"
    `include "json_number_test.svh"
    `include "json_array_test.svh"
    `include "json_object_test.svh"

    //`include "demo_test.svh"

endpackage

